`timescale 1ps/1ps

`include "header_systolic_2x2_2x2.sv"

// vcs -sverilog -full64 -timescale=1ns/1ps ../../../../../coredec_acc_soc/accelerator_soc/MeshMultiCgraRTL__explicit_systolic_2x2_2x2__pickled.v ../MeshMultiCgraRTL_systolic_2x2_2x2_tb.v -debug_access+all +incdir+..

module cgra_test
(
);

  logic [0:0] clk;
  logic [0:0] reset;

  IntraCgraPacket_4_2x2_4_8_2_CgraPayload__23265230afd8a14d recv_from_cpu_pkt__msg;
  logic [0:0] recv_from_cpu_pkt__rdy;
  logic [0:0] recv_from_cpu_pkt__val;

  IntraCgraPacket_4_2x2_4_8_2_CgraPayload__23265230afd8a14d send_to_cpu_pkt__msg;
  logic [0:0] send_to_cpu_pkt__rdy;
  logic [0:0] send_to_cpu_pkt__val;

  MeshMultiCgraRTL__explicit_systolic_2x2_2x2__pickled MultiCGRA (.*);

  int  PASS         = 'd0;
  time pass_time_of = 'd0;

  initial
  begin
    $display("\nTEST begin\n");

    clk = 1'b0;
    recv_from_cpu_pkt__val = 1'b0;
    send_to_cpu_pkt__rdy   = 1'b1;

    reset = 1'b0;
    #7
    reset = 1'b1;
    #50
    reset = 1'b0;
    #10
/*
typedef struct packed {
  logic [2:0] src;
  logic [2:0] dst;
  logic [1:0] src_cgra_id;
  logic [1:0] dst_cgra_id;
  logic [0:0] src_cgra_x;
  logic [0:0] src_cgra_y;
  logic [0:0] dst_cgra_x;
  logic [0:0] dst_cgra_y;
  logic [7:0] opaque;
  logic [0:0] vc_id;
  MultiCgraPayload_Cmd_Data_DataAddr_Ctrl_CtrlAddr__d9140faa89010e06 payload;
} IntraCgraPacket_4_2x2_4_8_2_CgraPayload__23265230afd8a14d;
*/
/*
typedef struct packed {
  logic [5:0] cmd;
  CgraData_32_1_1_1__payload_32__predicate_1__bypass_1__delay_1 data;
  logic [6:0] data_addr;
  CGRAConfig_7_4_2_4_4_3__49d22cda396bec88 ctrl;
  logic [3:0] ctrl_addr;
} MultiCgraPayload_Cmd_Data_DataAddr_Ctrl_CtrlAddr__d9140faa89010e06;
*/
/*
typedef struct packed {
  logic [31:0] payload;
  logic [0:0] predicate;
  logic [0:0] bypass;
  logic [0:0] delay;
} CgraData_32_1_1_1__payload_32__predicate_1__bypass_1__delay_1;
*/
/*
typedef struct packed {
  logic [6:0] operation;
  logic [3:0][2:0] fu_in;
  logic [7:0][2:0] routing_xbar_outport;
  logic [7:0][1:0] fu_xbar_outport;
  logic [2:0] vector_factor_power;
  logic [0:0] is_last_ctrl;
  logic [3:0][1:0] write_reg_from;
  logic [3:0][3:0] write_reg_idx;
  logic [3:0][0:0] read_reg_from;
  logic [3:0][3:0] read_reg_idx;
} CGRAConfig_7_4_2_4_4_3__49d22cda396bec88;
*/

/*
    input logic [180:0] inp_recv_from_cpu_pkt__msg,
    input logic [0:0] ref_recv_from_cpu_pkt__rdy,
    input logic [0:0] inp_recv_from_cpu_pkt__val,
    input logic [180:0] ref_send_to_cpu_pkt__msg,
    input logic [0:0] inp_send_to_cpu_pkt__rdy,
    input logic [0:0] ref_send_to_cpu_pkt__val,
*/
    #10
    recv_from_cpu_pkt__val = 1'b1;
    recv_from_cpu_pkt__msg = unpack_pkt('h0110001800000003200000000000000000000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0110001800000005208000000000000000000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0110001800000007210000000000000000000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0010001800000009218000000000000000000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h001000180000000b220000000000000000000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h001000180000000d228000000000000000000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h010000180000000f000000000000000000000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0100001800000011008000000000000000000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0100001800000013010000000000000000000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0110001a00000081000000000000000000000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0110001a00000083000000000000000000000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0110001a00000085000000000000000000000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0110001000000003000000000000000000000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0110000e00000007000000000000000000000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0110000600000000001c8d100000000400000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0110000000000000000000000000000000000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0010001a00000087000000000000000000000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0010001a00000089000000000000000000000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0010001a0000008b000000000000000000000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0010001000000003000000000000000000000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0010000e00000007000000000000000000000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0010000600000000001c8d100000000400000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0010000000000000000000000000000000000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0100001a00000001000000000000000000000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0100001a00000003000000000000000000000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0100001a00000005000000000000000000000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0100001000000003000000000000000000000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0100000e00000007000000000000000000000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0100000600000000001c8d100000000400000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0100000000000000000000000000000000000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0190001a00000005000000000000000000000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0190001000000003000000000000000000000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0190000e00000007000000000000000000000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0190000600000000001d8d100360000040000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0190000000000000000000000000000000000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0090001a00000009000000000000000000000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0090001000000003000000000000000000000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0090000e00000007000000000000000000000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0090000600000000001e8d104360000040000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0090000000000000000000000000000000000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0180001a0000000d000000000000000000000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0180001000000003000000000000000000000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0180000e00000007000000000000000000000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0180000600000000001e8d104360000040000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0180000000000000000000000000000000000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0080001a00000007000000000000000000000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0080001a00000009000000000000000000000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0080001a0000000b000000000000000000000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0080001000000003000000000000000000000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0080000e00000007000000000000000000000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0080000600000000003a8d100100000000000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0080000000000000000000000000000000000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0118001a00000011000000000000000000000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0118001000000003000000000000000000000000000000,'h1,'h1,'h0a42001c00000000000000000000000000000000000000,'h1,'h1);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0118000e00000007000000000000000000000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0118000600000000001d8d100360000040000000000000,'h0,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0118000600000000001d8d100360000040000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0118000000000000000000000000000000000000000000,'h1,'h1,'h0000000000000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0018001a00000015000000000000000000000000000000,'h1,'h1,'h0242001c00000000000000000000000000000000000000,'h1,'h1);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0018001000000003000000000000000000000000000000,'h0,'h1,'h0a00001c00000000000000000000000000000000000000,'h1,'h1);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0018001000000003000000000000000000000000000000,'h1,'h1,'h0242001c00000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0018000e00000007000000000000000000000000000000,'h1,'h1,'h0242001c00000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0018000600000000001e8d104360000040000000000000,'h1,'h1,'h0242001c00000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0018000000000000000000000000000000000000000000,'h1,'h1,'h0242001c00000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0108001a00000019000000000000000000000000000000,'h1,'h1,'h0242001c00000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0108001000000003000000000000000000000000000000,'h1,'h1,'h0242001c00000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0108000e00000007000000000000000000000000000000,'h1,'h1,'h0242001c00000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0108000600000000001e8d104360000040000000000000,'h1,'h1,'h0242001c00000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0108000000000000000000000000000000000000000000,'h1,'h1,'h0242001c00000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0008001a00000041000000000000000000000000000000,'h0,'h1,'h0600001c00000000000000000000000000000000000000,'h1,'h1);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0008001a00000041000000000000000000000000000000,'h1,'h1,'h0a00001c00000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0008001a00000043000000000000000000000000000000,'h1,'h1,'h0a00001c00000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0008001a00000045000000000000000000000000000000,'h1,'h1,'h0a00001c00000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0008001000000003000000000000000000000000000000,'h1,'h1,'h0a00001c00000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0008000e00000007000000000000000000000000000000,'h1,'h1,'h0a00001c00000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0008000600000000003a8d100100000000000000000000,'h1,'h1,'h0a00001c00000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0008000000000000000000000000000000000000000000,'h1,'h1,'h0a00001c00000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0198001a0000001d000000000000000000000000000000,'h1,'h1,'h0a00001c00000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0198001000000003000000000000000000000000000000,'h1,'h1,'h0a00001c00000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0198000e00000007000000000000000000000000000000,'h1,'h1,'h0e42001c00000000000000000000000000000000000000,'h1,'h1);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0198000600000000001d8d100300000040000000000000,'h1,'h1,'h0600001c00000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0198000000000000000000000000000000000000000000,'h1,'h1,'h0600001c00000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0098001a00000021000000000000000000000000000000,'h1,'h1,'h0600001c00000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0098001000000003000000000000000000000000000000,'h1,'h1,'h0600001c00000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0098000e00000007000000000000000000000000000000,'h1,'h1,'h0642001c00000000000000000000000000000000000000,'h1,'h1);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0098000600000000001e8d104300000040000000000000,'h1,'h1,'h0e42001c00000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0098000000000000000000000000000000000000000000,'h0,'h1,'h0e00001c00000000000000000000000000000000000000,'h1,'h1);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0098000000000000000000000000000000000000000000,'h1,'h1,'h0642001c00000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0188001a00000025000000000000000000000000000000,'h1,'h1,'h0642001c00000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0188001000000003000000000000000000000000000000,'h1,'h1,'h0642001c00000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0188000e00000007000000000000000000000000000000,'h1,'h1,'h0642001c00000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0188000600000000001e8d104300000040000000000000,'h1,'h1,'h0642001c00000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0188000000000000000000000000000000000000000000,'h1,'h1,'h0642001c00000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0088001a00000047000000000000000000000000000000,'h1,'h1,'h0642001c00000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0088001a00000049000000000000000000000000000000,'h1,'h1,'h0642001c00000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0088001a0000004b000000000000000000000000000000,'h1,'h1,'h0224001c00000000000000000000000000000000000000,'h1,'h1);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0088001000000003000000000000000000000000000000,'h1,'h1,'h0e00001c00000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0088000e00000007000000000000000000000000000000,'h1,'h1,'h0e00001c00000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0088000600000000003a8d100100000000000000000000,'h1,'h1,'h0e00001c00000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0088000000000000000000000000000000000000000000,'h1,'h1,'h0e00001c00000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0000001400000000018000000000000000000000000000,'h1,'h1,'h0e24001c00000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0000001400000000020000000000000000000000000000,'h1,'h1,'h0e24001c00000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0000001400000000028000000000000000000000000000,'h1,'h1,'h0e24001c00000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0000001400000000100000000000000000000000000000,'h1,'h1,'h0e24001c00000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0000001400000000108000000000000000000000000000,'h1,'h1,'h0e24001c00000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0000001400000000110000000000000000000000000000,'h1,'h1,'h0e24001c00000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0000001400000000118000000000000000000000000000,'h1,'h1,'h0e24001c00000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0000001400000000120000000000000000000000000000,'h0,'h1,'h0e24001c00000000000000000000000000000000000000,'h1,'h0);
    #10 // duplicate
    recv_from_cpu_pkt__msg = unpack_pkt('h0000001400000000120000000000000000000000000000,'h0,'h1,'h0e24001c00000000000000000000000000000000000000,'h1,'h0);
    #10 // triplicate
    recv_from_cpu_pkt__msg = unpack_pkt('h0000001400000000120000000000000000000000000000,'h1,'h1,'h0e24001c00000000000000000000000000000000000000,'h1,'h0);
    #10
    recv_from_cpu_pkt__msg = unpack_pkt('h0000001400000000128000000000000000000000000000,'h0,'h1,'h0200001600000079018000000000000000000000000000,'h1,'h1);
    #10 // duplicate
    recv_from_cpu_pkt__msg = unpack_pkt('h0000001400000000128000000000000000000000000000,'h1,'h1,'h0624001c00000000000000000000000000000000000000,'h1,'h0);
    
    #10
    recv_from_cpu_pkt__val = 0;

    #3000

    if ('d1 == PASS) $display("TEST PASSED at %0t.", pass_time_of);
    else             $display("TEST FAILED at %0t.", $time);

    $display("#########cgra 0 tile 0 cnst mem#################");
    for (int i = 0; i < 512; i++)
    begin
      if ( !$isunknown(MultiCGRA.cgra__0.tile__0.const_mem.reg_file.regs[i]) )
        $display("cgra0tile0cnst %d %d %d (%d)", i, MultiCGRA.cgra__0.tile__0.const_mem.reg_file.regs[i].payload, MultiCGRA.cgra__0.tile__0.const_mem.reg_file.regs[i].predicate, MultiCGRA.cgra__0.tile__0.const_mem.reg_file.regs[i]);
    end
    $display("##########################");
    for (int i = 0; i < 512; i++)
    begin
      if ( !$isunknown(MultiCGRA.cgra__0.tile__1.const_mem.reg_file.regs[i]) )
        $display("cgra0tile1cnst %d %d", i, MultiCGRA.cgra__0.tile__1.const_mem.reg_file.regs[i]);
    end
    $display("##########################");
    
    $display("********cgra 0 ctrl mem******************");
    for (int i = 0; i < 512; i++)
    begin
      if ( !$isunknown(MultiCGRA.cgra__0.tile__0.ctrl_mem.reg_file.regs[i]) )
        $display("cgra0tile0ctrl %d %d", i, MultiCGRA.cgra__0.tile__0.ctrl_mem.reg_file.regs[i]);
    end
    $display("##########################");
    for (int i = 0; i < 512; i++)
    begin
      if ( !$isunknown(MultiCGRA.cgra__0.tile__1.ctrl_mem.reg_file.regs[i]) )
        $display("cgra0tile1ctrl %d %d", i, MultiCGRA.cgra__0.tile__1.ctrl_mem.reg_file.regs[i]);
    end
    $display("##########################");
    
    $display("*************cgra0 data mem 0*************");
    for (int i = 0; i < 16; i++)
    begin
      if ( !$isunknown(MultiCGRA.cgra__0.data_mem.memory_wrapper__0.memory.regs[i]) )
        $display("cgra0regfile0 (addr 0 init) %d %d (%d)", i, MultiCGRA.cgra__0.data_mem.memory_wrapper__0.memory.regs[i].payload, MultiCGRA.cgra__0.data_mem.memory_wrapper__0.memory.regs[i]);
    end
    $display("#############cgra0 data mem 1#############");
    for (int i = 0; i < 16; i++)
    begin
      if ( !$isunknown(MultiCGRA.cgra__0.data_mem.memory_wrapper__1.memory.regs[i]) )
        $display("cgra0regfile1 (addr 0 init) %d %d", i, MultiCGRA.cgra__0.data_mem.memory_wrapper__1.memory.regs[i]);
    end

    $finish();
  end

  initial
    forever
    begin
      #5
      clk = ~clk;
    end

  always @ (posedge clk or negedge clk)
  begin
    #1

    if ( send_to_cpu_pkt__val && ('d300 == send_to_cpu_pkt__msg.payload.data.payload) && ('d1 == send_to_cpu_pkt__msg.payload.data.predicate) )
    begin
      PASS         = 'd1;
      pass_time_of = $time;
    end
  end

  /*initial
  begin  
    $dumpfile("./output.vcd");
    $dumpvars (0, cgra_test);
  end*/
  // The Verilator test fails on these $fsdb* functions; if pragmas do not work, add --bbox-sys to Verilator cmd.
`ifndef VERILATOR
  initial
  begin
    $fsdbDumpfile("./output.fsdb");
    $fsdbDumpvars ("+all", "cgra_test");
    $fsdbDumpMDA;
    $fsdbDumpSVA;
  end
`endif


endmodule

